--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY disp_rst IS PORT(clk:IN std_logic;rst_n:IN std_logic;done:OUT std_logic;s_rst:OUT std_logic);END disp_rst ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE fsm OF disp_rst IS SIGNAL z1b95a78d9:integer RANGE 1 DOWNTO 0;TYPE STATE_TYPE IS(z64ab6e507,zcc57584f0,zfdf6b4fa1,z6ecc89d31);SIGNAL zdf0be1ce6:STATE_TYPE;SIGNAL ze8e79043b:STATE_TYPE;SIGNAL zddc9dc0bc:std_logic_vector(6 DOWNTO 0);SIGNAL z28618b6b9:std_logic_vector(6 DOWNTO 0);SIGNAL za21ed1d6a:std_logic;SIGNAL z2e513ad1b:std_logic;SIGNAL zf3c003a58:std_logic;BEGIN z9149816e0:PROCESS(clk,rst_n)BEGIN IF(rst_n='0')THEN zdf0be1ce6<=z6ecc89d31;zddc9dc0bc<=(OTHERS=>'0');z1b95a78d9<=0;ELSIF(clk'EVENT AND clk='1')THEN zdf0be1ce6<=ze8e79043b;zddc9dc0bc<=z28618b6b9;CASE zdf0be1ce6 IS WHEN zcc57584f0=>z1b95a78d9<=1;WHEN OTHERS=>NULL;END CASE;END IF;END PROCESS z9149816e0;z145fbcc0d:PROCESS(za21ed1d6a,zdf0be1ce6,z1b95a78d9)BEGIN z2e513ad1b<='0';zf3c003a58<='0';CASE zdf0be1ce6 IS WHEN z64ab6e507=>IF(za21ed1d6a='1'AND(z1b95a78d9=1))THEN ze8e79043b<=zfdf6b4fa1;ELSIF(za21ed1d6a='1')THEN ze8e79043b<=zcc57584f0;zf3c003a58<='1';ELSE ze8e79043b<=z64ab6e507;END IF;WHEN zcc57584f0=>IF(za21ed1d6a='1')THEN ze8e79043b<=z64ab6e507;z2e513ad1b<='1';ELSE ze8e79043b<=zcc57584f0;END IF;WHEN zfdf6b4fa1=>ze8e79043b<=zfdf6b4fa1;WHEN z6ecc89d31=>ze8e79043b<=z64ab6e507;z2e513ad1b<='1';WHEN OTHERS=>ze8e79043b<=z6ecc89d31;END CASE;END PROCESS z145fbcc0d;z822bdb2c3:PROCESS(zdf0be1ce6)BEGIN done<='0';s_rst<='1';CASE zdf0be1ce6 IS WHEN z64ab6e507=>s_rst<='1';WHEN zcc57584f0=>s_rst<='0';WHEN zfdf6b4fa1=>done<='1';WHEN OTHERS=>NULL;END CASE;END PROCESS z822bdb2c3;zc4c7d2805:PROCESS(zddc9dc0bc,z2e513ad1b,zf3c003a58)VARIABLE z35e1a2c8c:std_logic;BEGIN IF(unsigned(zddc9dc0bc)=0)THEN z35e1a2c8c:='1';ELSE z35e1a2c8c:='0';END IF;IF(z2e513ad1b='1')THEN z28618b6b9<="1100011";ELSIF(zf3c003a58='1')THEN z28618b6b9<="1100011";ELSE IF(z35e1a2c8c='1')THEN z28618b6b9<=(OTHERS=>'0');ELSE z28618b6b9<=unsigned(zddc9dc0bc)-'1';END IF;END IF;za21ed1d6a<=z35e1a2c8c;END PROCESS zc4c7d2805;END fsm;