--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY disp_serial_led_cannon IS PORT(clk:IN std_logic;pixdata:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic;run:IN std_logic;bit_out:OUT std_logic;chans:OUT std_logic_vector(7 DOWNTO 0);lat:OUT std_logic;tx:OUT std_logic;y:OUT std_logic_vector(7 DOWNTO 0);x:OUT std_logic_vector(7 DOWNTO 0));END disp_serial_led_cannon ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE fsm OF disp_serial_led_cannon IS SIGNAL z1f2574037:std_logic_vector(7 DOWNTO 0);SIGNAL zbddb18e97:integer RANGE 23 DOWNTO-1;TYPE STATE_TYPE IS(z300f5740b,z82451b49a,z5b4a4026f,z40d04e6e4,z3638d9054,zd7d061bae,z8d5d87383,z6f19eeb13,zda3721a5d,z811b67cb9,zfed9561eb,z1b7cf85f1,zc42e36d33);SIGNAL zdf0be1ce6:STATE_TYPE;SIGNAL ze8e79043b:STATE_TYPE;SIGNAL zddc9dc0bc:std_logic_vector(12 DOWNTO 0);SIGNAL z28618b6b9:std_logic_vector(12 DOWNTO 0);SIGNAL za21ed1d6a:std_logic;SIGNAL z3f442e4ea:std_logic;SIGNAL z145d2d1b7:std_logic;SIGNAL z4fc46770e:std_logic;SIGNAL z4d1a0fb73:std_logic_vector(7 DOWNTO 0);SIGNAL z504ac3a28:std_logic_vector(7 DOWNTO 0);SIGNAL zdfaf1c3b8:std_logic_vector(7 DOWNTO 0);BEGIN z9149816e0:PROCESS(clk,rst_n)BEGIN IF(rst_n='0')THEN zdf0be1ce6<=z300f5740b;zddc9dc0bc<=(OTHERS=>'0');z4d1a0fb73<="00000000";z504ac3a28<="00000001";zdfaf1c3b8<="00000001";z1f2574037<="00000000";zbddb18e97<=23;ELSIF(clk'EVENT AND clk='1')THEN zdf0be1ce6<=ze8e79043b;zddc9dc0bc<=z28618b6b9;CASE zdf0be1ce6 IS WHEN z5b4a4026f=>zbddb18e97<=zbddb18e97-1;WHEN zd7d061bae=>z504ac3a28<=z504ac3a28(6 downto 0)&'0';zbddb18e97<=23;WHEN z8d5d87383=>zdfaf1c3b8<=zdfaf1c3b8(6 downto 0)&'0';z504ac3a28<="00000001";zbddb18e97<=23;WHEN z6f19eeb13=>z1f2574037<=z1f2574037(6 downto 0)&'0';WHEN zda3721a5d=>z504ac3a28<="00000001";zdfaf1c3b8<="00000001";zbddb18e97<=23;WHEN z811b67cb9=>z1f2574037<="00000001";WHEN z1b7cf85f1=>z4d1a0fb73<=z1f2574037;WHEN zc42e36d33=>z4d1a0fb73<="00000000";WHEN OTHERS=>NULL;END CASE;END IF;END PROCESS z9149816e0;z145fbcc0d:PROCESS(z1f2574037,za21ed1d6a,zdf0be1ce6,zbddb18e97,run,z504ac3a28,zdfaf1c3b8)BEGIN z3f442e4ea<='0';z145d2d1b7<='0';z4fc46770e<='0';CASE zdf0be1ce6 IS WHEN z300f5740b=>IF(run='1')THEN ze8e79043b<=z82451b49a;ELSE ze8e79043b<=z300f5740b;END IF;WHEN z82451b49a=>IF(run='0')THEN ze8e79043b<=z5b4a4026f;ELSE ze8e79043b<=z82451b49a;END IF;WHEN z5b4a4026f=>ze8e79043b<=z3638d9054;WHEN z40d04e6e4=>IF(za21ed1d6a='1')THEN ze8e79043b<=z6f19eeb13;ELSE ze8e79043b<=z40d04e6e4;END IF;WHEN z3638d9054=>IF(z504ac3a28="10000000"AND zdfaf1c3b8="10000000"AND zbddb18e97=-1)THEN ze8e79043b<=zda3721a5d;ELSIF(z504ac3a28="10000000"AND zbddb18e97=-1)THEN ze8e79043b<=z8d5d87383;ELSIF(zbddb18e97=-1)THEN ze8e79043b<=zd7d061bae;ELSE ze8e79043b<=z300f5740b;END IF;WHEN zd7d061bae=>ze8e79043b<=z300f5740b;WHEN z8d5d87383=>ze8e79043b<=zc42e36d33;z4fc46770e<='1';WHEN z6f19eeb13=>ze8e79043b<=zfed9561eb;WHEN zda3721a5d=>ze8e79043b<=zc42e36d33;z4fc46770e<='1';WHEN z811b67cb9=>ze8e79043b<=z1b7cf85f1;z145d2d1b7<='1';WHEN zfed9561eb=>IF(z1f2574037="00000000")THEN ze8e79043b<=z811b67cb9;ELSE ze8e79043b<=z1b7cf85f1;z145d2d1b7<='1';END IF;WHEN z1b7cf85f1=>ze8e79043b<=z300f5740b;WHEN zc42e36d33=>IF(za21ed1d6a='1')THEN ze8e79043b<=z40d04e6e4;z3f442e4ea<='1';ELSE ze8e79043b<=zc42e36d33;END IF;WHEN OTHERS=>ze8e79043b<=z300f5740b;END CASE;END PROCESS z145fbcc0d;z822bdb2c3:PROCESS(zdf0be1ce6,zbddb18e97,pixdata)BEGIN bit_out<='0';lat<='0';tx<='0';CASE zdf0be1ce6 IS WHEN z82451b49a=>bit_out<=pixdata(zbddb18e97);tx<='1';WHEN z40d04e6e4=>lat<='1';WHEN OTHERS=>NULL;END CASE;END PROCESS z822bdb2c3;zc4c7d2805:PROCESS(zddc9dc0bc,z3f442e4ea,z145d2d1b7,z4fc46770e)VARIABLE z35e1a2c8c:std_logic;BEGIN IF(unsigned(zddc9dc0bc)=0)THEN z35e1a2c8c:='1';ELSE z35e1a2c8c:='0';END IF;IF(z3f442e4ea='1')THEN z28618b6b9<="0000000000011";ELSIF(z145d2d1b7='1')THEN z28618b6b9<="1011000100001";ELSIF(z4fc46770e='1')THEN z28618b6b9<="0111110011111";ELSE IF(z35e1a2c8c='1')THEN z28618b6b9<=(OTHERS=>'0');ELSE z28618b6b9<=unsigned(zddc9dc0bc)-'1';END IF;END IF;za21ed1d6a<=z35e1a2c8c;END PROCESS zc4c7d2805;chans<=z4d1a0fb73;y<=z504ac3a28;x<=zdfaf1c3b8;END fsm;